`define SIMULATION
// `define NOCACHE
// `define DISABLE_PIPELINE


// Uncomment to use this configuration, ONLY 1 AT A TIME!!!
`define SINGLECORE
// `define MULTICORE2
// `define MULTICORE4