module vfm_proc_inst(
    input [1:0] push_button,
    input [3:0] dip_switchs,
    output reg LEDS

);



endmodule